module entradas ( 
	a,
	b,
	c,
	d,
	e,
	f1,
	f2,
	f3,
	f4,
	f5,
	f6
	) ;

input  a;
input  b;
input  c;
input  d;
input  e;
inout  f1;
inout  f2;
inout  f3;
inout  f4;
inout  f5;
inout  f6;
