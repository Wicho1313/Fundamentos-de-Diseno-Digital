module deco ( 
	e,
	display
	) ;

input [2:0] e;
inout [6:0] display;
