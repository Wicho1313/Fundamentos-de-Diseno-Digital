module aritmeticos ( 
	a,
	b,
	c,
	semisuma,
	suma,
	semiresta,
	resta,
	multi,
	c1,
	c2,
	c3,
	c4
	) ;

input  a;
input  b;
input  c;
inout  semisuma;
inout  suma;
inout  semiresta;
inout  resta;
inout  multi;
inout  c1;
inout  c2;
inout  c3;
inout  c4;
