LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ARITMETICOS IS
	PORT(A, B, C: IN STD_LOGIC; 
	SEMISUMA, SUMA, SEMIRESTA, RESTA, MULTI, C1, C2, C3, C4: OUT STD_LOGIC);
END ARITMETICOS;

ARCHITECTURE CIRCUITOS OF ARITMETICOS IS
BEGIN
	SEMISUMA <= A XOR B;
	C1 <= A AND B;
	SUMA <= A XOR B XOR C;
	C2 <= (A AND B) OR (B AND C) OR (A AND C);
	SEMIRESTA <= A XOR B;
	C3 <= (NOT A) AND B;
	RESTA <= A XOR B XOR C;
	C4 <= ((NOT A) AND B) OR (B AND C) OR ((NOT A) AND C);
END CIRCUITOS;


